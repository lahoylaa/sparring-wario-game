
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package package_end_pos_2 is
    constant IMAGE_WIDTH  : integer := 50;
    constant IMAGE_HEIGHT : integer := 50;
    type image_array is array (0 to 2499) of std_logic_vector(15 downto 0);
    constant end_pos_2 : image_array := (
   "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111001110001010",
        "1111111111111111",
        "1111001110001010",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111111111110000",
        "1111111111111111",
        "1111111111111111",
        "1111111111110000",
        "1111101110110000",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111001110001010",
        "1111111111111111",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111010100010000",
        "1111111111111111",
        "1111001110001010",
        "1111001110001010",
        "1111000000000000",
        "1111111111111111",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111010100010000",
        "1111101110110000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111010100010000",
        "1111111111111111",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111010100010000",
        "1111101110111011",
        "1111010100010000",
        "1111010100010000",
        "1111101110111011",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111101110110000",
        "1111111111110000",
        "1111111111110000",
        "1111010100010000",
        "1111111111111111",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111101110110000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111111111110000",
        "1111101110110000",
        "1111010100010000",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111010100010000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111010100010000",
        "1111001110001010",
        "1111001110001010",
        "1111010100010000",
        "1111000100001101",
        "1111111111110000",
        "1111101100000000",
        "1111000100001101",
        "1111101100000000",
        "1111111111110000",
        "1111000100001101",
        "1111101110110000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110110000",
        "1111010100010000",
        "1111010100010000",
        "1111101100000000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111010100010000",
        "1111010100010000",
        "1111101110110000",
        "1111111111110000",
        "1111000100001101",
        "1111101100000000",
        "1111000100001101",
        "1111101100000000",
        "1111000100001101",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111101110110000",
        "1111010100010000",
        "1111101100000000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000100001101",
        "1111101100000000",
        "1111000100001101",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111111111111111",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110111011",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111101110111011",
        "1111101110000110",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101100000000",
        "1111111100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "1111001110001010",
        "1111101110111011",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111111111111111",
        "1111101110111011",
        "1111101110111011",
        "1111001110001010",
        "1111101110000110",
        "1111101100000000",
        "1111111100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111010010101110",
        "1111111111111111",
        "1111000000000000",
        "1111111111111111",
        "1111000000000000",
        "1111101110000110",
        "1111000000000000",
        "1111101110111011",
        "1111111111111111",
        "1111000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111010010101110",
        "1111101110000110",
        "1111101100000000",
        "1111111100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111001110001010",
        "1111111111111111",
        "1111111111111111",
        "1111101110111011",
        "1111000000000000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110111011",
        "1111111111111111",
        "1111111111111111",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111101100000000",
        "1111111100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111111010010111",
        "1111101110000110",
        "1111010010101110",
        "1111111010010111",
        "1111010100010000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111111100000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111111010010111",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111101100000000",
        "1111111101111011",
        "1111111100000000",
        "1111111100000000",
        "1111111100000000",
        "1111101100000000",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111111100000000",
        "1111010100010000",
        "1111101110110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111010100010000",
        "1111101100000000",
        "1111111101111011",
        "1111111111111111",
        "1111111101111011",
        "1111111100000000",
        "1111111100000000",
        "1111111100000000",
        "1111101100000000",
        "1111010100010000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111101110110000",
        "1111111111110000",
        "1111111111111111",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111101100000000",
        "1111101100000000",
        "1111111101111011",
        "1111111100000000",
        "1111111100000000",
        "1111111100000000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111000000000000",
        "1111010100010000",
        "1111101110110000",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111101100000000",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101110110000",
        "1111111111111111",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101110110000",
        "1111101110110000",
        "1111111111110000",
        "1111111111110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111000000000000",
        "1111101110000110",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111111111111111",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111010100010000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111111010010111",
        "1111010100010000",
        "1111000000000000",
        "1111101110111011",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111101110110000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000000000",
        "1111111010010111",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111111111111111",
        "1111111111111111",
        "1111101110111011",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111101110111011",
        "1111000000000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111010100010000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110111011",
        "1111101110111011",
        "1111000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111101110111011",
        "1111000000000000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111010010101110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000000000",
        "1111111010010111",
        "1111111010010111",
        "1111010100010000",
        "1111101110111011",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111101110111011",
        "1111111111111111",
        "1111101110111011",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111010010111",
        "1111010100010000",
        "1111000000000000",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111101110111011",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010010101110",
        "1111010100010000",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111111010010111",
        "1111111010010111",
        "1111101110000110",
        "1111010100010000",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111000000001001",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111111010010111",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111111010010111",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111111010010111",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111010010101110",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111001110001010",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111001110001010",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111001110001010",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111001110001010",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111001110001010",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111010100010000",
        "1111001110001010",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111010010101110",
        "1111001110001010",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111001110001010",
        "1111001110001010",
        "1111010100010000",
        "1111001110001010",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111010010101110",
        "1111001110001010",
        "1111001110001010",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111010100010000",
        "1111001110001010",
        "1111001110001010",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111010010101110",
        "1111001110001010",
        "1111001110001010",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111001110001010",
        "1111010100010000",
        "1111001110001010",
        "1111001110001010",
        "1111001110001010",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111101110000110",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111101110000110",
        "1111010100010000",
        "1111010100010000",
        "1111010100010000",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111111101111011",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111010100010000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000001001",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111111101111011",
        "1111101110000110",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111101110000110",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000001001",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "1111000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000"
    );
end package package_end_pos_2;