library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package package_ball_pink is
    constant IMAGE_WIDTH  : integer := 20;
    constant IMAGE_HEIGHT : integer := 20;
    type image_array is array (0 to 399) of std_logic_vector(15 downto 0);
    constant ball_pink : image_array := (
          "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111100000101",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111101111001",
        "1111111110101100",
        "1111111110101100",
        "1111111110101100",
        "1111111110101100",
        "1111111110101100",
        "1111111110101100",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111110101100",
        "1111111111101110",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111110101100",
        "1111111111101110",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111110101100",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111101111001",
        "1111111111101110",
        "1111111110101100",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111100000101",
        "1111111100000101",
        "1111111101111001",
        "1111111101111001",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111100000101",
        "1111111111111111",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "1111111111111111",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000",
        "0000000000000000"
    );
end package package_ball_pink;